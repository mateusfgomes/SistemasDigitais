CASE estado IS
						WHEN cents100 =>
							estado <= refri;
							display_2 <= "1000000"; -- 0
							display_1 <= "1000000"; -- 0
							display_0 <= "1000000";	-- 0
						WHEN cents95 =>
							estado <= cents0;
							display_0 <= "1000000";	-- 0
							display_1 <= "0010000"; -- 9
							display_2 <= "0010010"; -- 5
						WHEN cents90 =>
							estado <= cents0;
							display_0 <= "1000000";	-- 0
							display_1 <= "0010000"; -- 9
							display_2 <= "1000000";	-- 0
						WHEN cents85 =>
							estado <= cents0;
							display_0 <= "1000000";	-- 0
							display_1 <= "0000000"; -- 8
							display_2 <= "0010010"; -- 5
						WHEN cents80 =>
							estado <= cents0;
							display_0 <= "1000000";	-- 0
							display_1 <= "0000000"; -- 8 
							display_2 <= "1000000";	-- 0
						WHEN cents75 =>
							estado <= cents0;
							display_0 <= "1000000";	-- 0
							display_1 <= "1111000"; -- 7
							display_1 <= "0010010"; -- 5
						WHEN cents70 =>
							estado <= cents0;
							display_0 <= "1000000";	-- 0
							display_1 <= "1111000"; -- 7
							display_2 <= "1000000";	-- 0
						WHEN cents65 =>
							estado <= cents0;
							display_0 <= "1000000";	-- 0
							display_1 <= "0000010"; -- 6
							display_2 <= "0010010"; -- 5
						WHEN cents60 =>
							estado <= cents0;
							display_0 <= "1000000";	-- 0
							display_1 <= "0000010"; -- 6
							display_2 <= "1000000";	-- 0
						WHEN cents55 =>
							estado <= cents0;
							display_0 <= "1000000";	-- 0
							display_1 <= "0010010"; -- 5
							display_2 <= "0010010"; -- 5
						WHEN cents50 =>
							estado <= cents0;
							display_0 <= "1000000";	-- 0
							display_1 <= "0010010"; -- 5
							display_2 <= "1000000";	-- 0
						WHEN cents45 =>
							estado <= cents0;
							display_0 <= "1000000";	-- 0
							display_1 <= "0011001"; -- 4
							display_2 <= "0010010"; -- 5
						WHEN cents40 =>
							estado <= cents0;
							display_0 <= "1000000";	-- 0
							display_1 <= "0011001"; -- 4
							display_2 <= "1000000";	-- 0
						WHEN cents35 =>
							estado <= cents0;
							display_0 <= "1000000";	-- 0
							display_1 <= "0110000"; -- 3
							display_2 <= "0010010"; -- 5
						WHEN cents30 =>
							estado <= cents0;
							display_0 <= "1000000";	-- 0
							display_1 <= "0110000"; -- 3
							display_2 <= "1000000";	-- 0
						WHEN cents25 =>
							estado <= cents0;
							display_0 <= "1000000";	-- 0
							display_1 <= "0100100"; -- 2
							display_2 <= "0010010"; -- 5
						WHEN cents20 =>
							estado <= cents0;
							display_0 <= "1000000";	-- 0
							display_1 <= "0100100"; -- 2
							display_2 <= "1000000";	-- 0
						WHEN cents10 =>
							estado <= cents0;
							display_0 <= "1000000";	-- 0
							display_1 <= "1111001"; -- 1
							display_2 <= "1000000";	-- 0
						WHEN cents0 =>
							estado <= cents0;
							display_0 <= "1000000";	-- 0
							display_1 <= "1000000";	-- 0
							display_2 <= "1000000";	-- 0
						WHEN refri =>
							estado <= refri;
							display_0 <= "1000000";	-- 0
							display_1 <= "1000000";	-- 0
							display_2 <= "1000000";	-- 0
					END CASE;